class BusOp;
	typedef enum {BYTE,WORD,LWRD} length_e;
	rand length_e len;
	