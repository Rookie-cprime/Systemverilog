library verilog;
use verilog.vl_types.all;
entity fetch_ifc is
    port(
        clk             : in     vl_logic
    );
end fetch_ifc;
