library verilog;
use verilog.vl_types.all;
entity test_1 is
end test_1;
