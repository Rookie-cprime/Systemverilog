/*************************************************
void和null类型的值和您在C语言中找到的值相同，void在函数中不返回值。
其中as null用于将变量与空值进行比较，例如将字符串与空字符串进行比较。
我们将在探索类数据类型时讨论这个问题。

chandle数据类型用于存储指针，同时使用直接编程接口。
我们将在DPI一节讨论这个问题。
**************************************************/