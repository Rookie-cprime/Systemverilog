library verilog;
use verilog.vl_types.all;
entity fetch_ifc_sv_unit is
end fetch_ifc_sv_unit;
